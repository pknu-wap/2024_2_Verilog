library verilog;
use verilog.vl_types.all;
entity tb_Cnt is
end tb_Cnt;
