library verilog;
use verilog.vl_types.all;
entity tb_Add4b is
end tb_Add4b;
