library verilog;
use verilog.vl_types.all;
entity tb_Add16b is
end tb_Add16b;
