library verilog;
use verilog.vl_types.all;
entity tb_AddSub4b is
end tb_AddSub4b;
