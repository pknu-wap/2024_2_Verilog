library verilog;
use verilog.vl_types.all;
entity tb_AddSub16b is
end tb_AddSub16b;
